`ifndef DSP
`define DSP

`define DSP_A 27
`define DSP_B 18
`define DSP_C 48
`define DSP_P 48

`define DSP_A_U (`DSP_A - 1)
`define DSP_B_U (`DSP_B - 1)
`define DSP_C_U (`DSP_C - 1)
`define DSP_M_U (`DSP_A_U + `DSP_B_U)

`endif