localparam DSP_A = 27,
localparam DSP_B = 18,
localparam DSP_C = 48,
localparam DSP_P = 48,


localparam DSP_A_U = DSP_A - 1,
localparam DSP_B_U = DSP_B - 1,
localparam DSP_C_U = DSP_C - 1,
localparam DSP_M_U = DSP_A_U + DSP_B_U
